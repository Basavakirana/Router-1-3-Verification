package router_test_pkg;

        // import the UVM package
        import uvm_pkg::*;

        // include the uvm_macros.svh
        `include "uvm_macros.svh"
        // include the tb_defs.sv
//        `include "tb_defs.sv"

        `include "source_transaction.sv"
        `include "source_agt_config.sv"
        `include "dest_agt_config.sv"
        `include "env_config.sv"
        `include "source_driver.sv"
        `include "source_monitor.sv"
        `include "source_sequencer.sv"
        `include "source_agt.sv"
        `include "source_agt_top.sv"
        `include "source_sequence.sv"

        `include "dest_transaction.sv"
        `include "dest_monitor.sv"
        `include "dest_sequencer.sv"
        `include "dest_sequence.sv"
        `include "dest_driver.sv"
        `include "dest_agt.sv"
        `include "dest_agt_top.sv"

        `include "router_vseqr.sv"
        `include "router_vseq.sv"
        `include "router_sb.sv"

        `include "router_env.sv"
        `include "router_test.sv"
endpackage
